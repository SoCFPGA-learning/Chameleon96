// soc_hps.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module soc_hps (
		output wire        clock_bridge_0_out_clk_clk,       // clock_bridge_0_out_clk.clk
		output wire [66:0] hps_0_h2f_loan_io_in,             //      hps_0_h2f_loan_io.in
		input  wire [66:0] hps_0_h2f_loan_io_out,            //                       .out
		input  wire [66:0] hps_0_h2f_loan_io_oe,             //                       .oe
		inout  wire        hps_io_hps_io_sdio_inst_CMD,      //                 hps_io.hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,       //                       .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,       //                       .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,      //                       .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,       //                       .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,       //                       .hps_io_sdio_inst_D3
		input  wire        hps_io_hps_io_uart0_inst_RX,      //                       .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,      //                       .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO14, //                       .hps_io_gpio_inst_LOANIO14
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO17, //                       .hps_io_gpio_inst_LOANIO17
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO19, //                       .hps_io_gpio_inst_LOANIO19
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO22, //                       .hps_io_gpio_inst_LOANIO22
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO23, //                       .hps_io_gpio_inst_LOANIO23
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO25, //                       .hps_io_gpio_inst_LOANIO25
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO27, //                       .hps_io_gpio_inst_LOANIO27
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO28, //                       .hps_io_gpio_inst_LOANIO28
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO29, //                       .hps_io_gpio_inst_LOANIO29
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO30, //                       .hps_io_gpio_inst_LOANIO30
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO32, //                       .hps_io_gpio_inst_LOANIO32
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO33, //                       .hps_io_gpio_inst_LOANIO33
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO34, //                       .hps_io_gpio_inst_LOANIO34
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO48, //                       .hps_io_gpio_inst_LOANIO48
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO53, //                       .hps_io_gpio_inst_LOANIO53
		inout  wire        hps_io_hps_io_gpio_inst_LOANIO54, //                       .hps_io_gpio_inst_LOANIO54
		output wire [14:0] memory_mem_a,                     //                 memory.mem_a
		output wire [2:0]  memory_mem_ba,                    //                       .mem_ba
		output wire        memory_mem_ck,                    //                       .mem_ck
		output wire        memory_mem_ck_n,                  //                       .mem_ck_n
		output wire        memory_mem_cke,                   //                       .mem_cke
		output wire        memory_mem_cs_n,                  //                       .mem_cs_n
		output wire        memory_mem_ras_n,                 //                       .mem_ras_n
		output wire        memory_mem_cas_n,                 //                       .mem_cas_n
		output wire        memory_mem_we_n,                  //                       .mem_we_n
		output wire        memory_mem_reset_n,               //                       .mem_reset_n
		inout  wire [15:0] memory_mem_dq,                    //                       .mem_dq
		inout  wire [1:0]  memory_mem_dqs,                   //                       .mem_dqs
		inout  wire [1:0]  memory_mem_dqs_n,                 //                       .mem_dqs_n
		output wire        memory_mem_odt,                   //                       .mem_odt
		output wire [1:0]  memory_mem_dm,                    //                       .mem_dm
		input  wire        memory_oct_rzqin                  //                       .oct_rzqin
	);

	soc_hps_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (0)
	) hps_0 (
		.h2f_loan_in               (hps_0_h2f_loan_io_in),             //     h2f_loan_io.in
		.h2f_loan_out              (hps_0_h2f_loan_io_out),            //                .out
		.h2f_loan_oe               (hps_0_h2f_loan_io_oe),             //                .oe
		.h2f_user0_clk             (clock_bridge_0_out_clk_clk),       // h2f_user0_clock.clk
		.mem_a                     (memory_mem_a),                     //          memory.mem_a
		.mem_ba                    (memory_mem_ba),                    //                .mem_ba
		.mem_ck                    (memory_mem_ck),                    //                .mem_ck
		.mem_ck_n                  (memory_mem_ck_n),                  //                .mem_ck_n
		.mem_cke                   (memory_mem_cke),                   //                .mem_cke
		.mem_cs_n                  (memory_mem_cs_n),                  //                .mem_cs_n
		.mem_ras_n                 (memory_mem_ras_n),                 //                .mem_ras_n
		.mem_cas_n                 (memory_mem_cas_n),                 //                .mem_cas_n
		.mem_we_n                  (memory_mem_we_n),                  //                .mem_we_n
		.mem_reset_n               (memory_mem_reset_n),               //                .mem_reset_n
		.mem_dq                    (memory_mem_dq),                    //                .mem_dq
		.mem_dqs                   (memory_mem_dqs),                   //                .mem_dqs
		.mem_dqs_n                 (memory_mem_dqs_n),                 //                .mem_dqs_n
		.mem_odt                   (memory_mem_odt),                   //                .mem_odt
		.mem_dm                    (memory_mem_dm),                    //                .mem_dm
		.oct_rzqin                 (memory_oct_rzqin),                 //                .oct_rzqin
		.hps_io_sdio_inst_CMD      (hps_io_hps_io_sdio_inst_CMD),      //          hps_io.hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0       (hps_io_hps_io_sdio_inst_D0),       //                .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1       (hps_io_hps_io_sdio_inst_D1),       //                .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK      (hps_io_hps_io_sdio_inst_CLK),      //                .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2       (hps_io_hps_io_sdio_inst_D2),       //                .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3       (hps_io_hps_io_sdio_inst_D3),       //                .hps_io_sdio_inst_D3
		.hps_io_uart0_inst_RX      (hps_io_hps_io_uart0_inst_RX),      //                .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX      (hps_io_hps_io_uart0_inst_TX),      //                .hps_io_uart0_inst_TX
		.hps_io_gpio_inst_LOANIO14 (hps_io_hps_io_gpio_inst_LOANIO14), //                .hps_io_gpio_inst_LOANIO14
		.hps_io_gpio_inst_LOANIO17 (hps_io_hps_io_gpio_inst_LOANIO17), //                .hps_io_gpio_inst_LOANIO17
		.hps_io_gpio_inst_LOANIO19 (hps_io_hps_io_gpio_inst_LOANIO19), //                .hps_io_gpio_inst_LOANIO19
		.hps_io_gpio_inst_LOANIO22 (hps_io_hps_io_gpio_inst_LOANIO22), //                .hps_io_gpio_inst_LOANIO22
		.hps_io_gpio_inst_LOANIO23 (hps_io_hps_io_gpio_inst_LOANIO23), //                .hps_io_gpio_inst_LOANIO23
		.hps_io_gpio_inst_LOANIO25 (hps_io_hps_io_gpio_inst_LOANIO25), //                .hps_io_gpio_inst_LOANIO25
		.hps_io_gpio_inst_LOANIO27 (hps_io_hps_io_gpio_inst_LOANIO27), //                .hps_io_gpio_inst_LOANIO27
		.hps_io_gpio_inst_LOANIO28 (hps_io_hps_io_gpio_inst_LOANIO28), //                .hps_io_gpio_inst_LOANIO28
		.hps_io_gpio_inst_LOANIO29 (hps_io_hps_io_gpio_inst_LOANIO29), //                .hps_io_gpio_inst_LOANIO29
		.hps_io_gpio_inst_LOANIO30 (hps_io_hps_io_gpio_inst_LOANIO30), //                .hps_io_gpio_inst_LOANIO30
		.hps_io_gpio_inst_LOANIO32 (hps_io_hps_io_gpio_inst_LOANIO32), //                .hps_io_gpio_inst_LOANIO32
		.hps_io_gpio_inst_LOANIO33 (hps_io_hps_io_gpio_inst_LOANIO33), //                .hps_io_gpio_inst_LOANIO33
		.hps_io_gpio_inst_LOANIO34 (hps_io_hps_io_gpio_inst_LOANIO34), //                .hps_io_gpio_inst_LOANIO34
		.hps_io_gpio_inst_LOANIO48 (hps_io_hps_io_gpio_inst_LOANIO48), //                .hps_io_gpio_inst_LOANIO48
		.hps_io_gpio_inst_LOANIO53 (hps_io_hps_io_gpio_inst_LOANIO53), //                .hps_io_gpio_inst_LOANIO53
		.hps_io_gpio_inst_LOANIO54 (hps_io_hps_io_gpio_inst_LOANIO54), //                .hps_io_gpio_inst_LOANIO54
		.h2f_rst_n                 ()                                  //       h2f_reset.reset_n
	);

endmodule
