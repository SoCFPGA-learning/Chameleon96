
module iOSC (
	oscena,
	clkout);	

	input		oscena;
	output		clkout;
endmodule
